module net

import time

const (
	no_deadline = time.Time{unix: 0}
)

pub struct TcpConn {
pub:
	sock TcpSocket

mut:
	write_deadline time.Time
	read_deadline time.Time

	read_timeout time.Duration
	write_timeout time.Duration
}

pub fn dial_tcp(address string) ?TcpConn {
	s := new_tcp_socket()?
	s.connect(address)?

	return TcpConn {
		sock: s
		
		read_timeout: -1
		write_timeout: -1
	}
}

pub fn (c TcpConn) close() ? {
	c.sock.close()?
	return none
}

// write blocks and attempts to write all data
pub fn (c TcpConn) write(bytes []byte) ? {
	unsafe {
		mut ptr_base := byteptr(bytes.data)
		mut total_sent := 0

		for total_sent < bytes.len {
			ptr := ptr_base + total_sent
			remaining := bytes.len - total_sent
			mut sent := C.send(c.sock.handle, ptr, remaining, msg_nosignal)

			if sent < 0 {
				code := error_code()
				match code {
					error_ewouldblock {
						c.wait_for_write()
						continue
					}
					else {
						wrap_error(code)?
					}
				}
			}
			total_sent += sent
		}
	}
	return none
}

pub fn (c TcpConn) read_into(mut buf []byte) ?int {
	res := C.recv(c.sock.handle, buf.data, buf.len, 0)

	if res >= 0 {
		return res
	}

	code := error_code()
	match code {
		error_ewouldblock {
			c.wait_for_read()?
			return socket_error(C.recv(c.sock.handle, buf.data, buf.len, 0))
		}
		else {
			wrap_error(code)?
		}
	}
}

pub fn (c TcpConn) read() ?[]byte {
	buf := []byte { len: 1024 }
	read := c.read_into(buf)?
	return buf[..read]
}

pub fn (c TcpConn) read_deadline() ?time.Time {
	if c.read_deadline.unix == 0 {
		return c.read_deadline
	}
	return none
}

pub fn (mut c TcpConn) set_read_deadline(deadline time.Time) {
	c.read_deadline = deadline
}

pub fn (c TcpConn) write_deadline() ?time.Time {
	if c.write_deadline.unix == 0 {
		return c.write_deadline
	}
	return none
}

pub fn (mut c TcpConn) set_write_deadline(deadline time.Time) {
	c.write_deadline = deadline
}

pub fn (c TcpConn) read_timeout() time.Duration {
	return c.read_timeout
}

pub fn(mut c TcpConn) set_read_timeout(t time.Duration) {
	c.read_timeout = t
}

pub fn (c TcpConn) write_timeout() time.Duration {
	return c.write_timeout
}

pub fn (mut c TcpConn) set_write_timeout(t time.Duration) {
	c.write_timeout = t
}

[inline]
pub fn (c TcpConn) wait_for_read() ? {
	return wait_for_read(c.sock.handle, c.read_deadline, c.read_timeout)
}

[inline]
pub fn (c TcpConn) wait_for_write() ? {
	return wait_for_write(c.sock.handle, c.write_deadline, c.write_timeout)
}

pub fn (c TcpConn) str() string {
	return ''
}

pub struct TcpListener {
	sock TcpSocket

mut:
	accept_timeout time.Duration
	accept_deadline time.Time
}

pub fn listen_tcp(port int) ?TcpListener {
	s := new_tcp_socket()?
	if port >= socket_max_port {
		return err_invalid_port
	}

	mut addr := C.sockaddr_in{}
	addr.sin_family = SocketFamily.inet
	addr.sin_port = C.htons(port)
	addr.sin_addr.s_addr = C.htonl(C.INADDR_ANY)
	size := sizeof(C.sockaddr_in)

	// cast to the correct type
	sockaddr := &C.sockaddr(&addr)

	socket_error(C.bind(s.handle, sockaddr, size))?
	socket_error(C.listen(s.handle, 128))?

	return TcpListener {
		sock: s
		accept_timeout: -1
		accept_deadline: no_deadline
	}
}

pub fn (l TcpListener) accept() ?TcpConn {
	addr := C.sockaddr_storage{}
	unsafe {
		C.memset(&addr, 0, sizeof(C.sockaddr_storage))
	}
	size := sizeof(C.sockaddr_storage)

	// cast to correct type
	sock_addr := &C.sockaddr(&addr)
	mut new_handle := C.accept(l.sock.handle, sock_addr, &size)

	if new_handle <= 0 {
		l.wait_for_accept()?

		new_handle = C.accept(l.sock.handle, sock_addr, &size)
		
		if new_handle == -1 || new_handle == 0 {
			return none
		}
	}

	new_sock := TcpSocket {
		handle: new_handle
	}

	return TcpConn{
		sock: new_sock
		read_timeout: -1
		write_timeout: -1
	}
}

pub fn (c TcpListener) accept_deadline() ?time.Time {
	if c.accept_deadline.unix != 0 {
		return c.accept_deadline
	}
	return none
}

pub fn (mut c TcpListener) set_accept_deadline(deadline time.Time) {
	c.accept_deadline = deadline
}

pub fn (c TcpListener) accept_timeout() time.Duration {
	return c.accept_timeout
}

pub fn(mut c TcpListener) set_accept_timeout(t time.Duration) {
	c.accept_timeout = t
}

pub fn (c TcpListener) wait_for_accept() ? {
	return wait_for_read(c.sock.handle, c.accept_deadline, c.accept_timeout)
}

pub fn (c TcpListener) close() ? {
	c.sock.close()?
	return none
}

struct TcpSocket {
pub:
	handle int
}

fn new_tcp_socket() ?TcpSocket {
	sockfd := socket_error(C.socket(SocketFamily.inet, SocketType.tcp, 0))?
	s := TcpSocket {
		handle: sockfd
	}
	s.set_option_bool(.reuse_addr, true)?
	$if windows {
		t := true
		socket_error(C.ioctlsocket(sockfd, fionbio, &t))?
	} $else {
		socket_error(C.fcntl(sockfd, C.F_SETFD, C.O_NONBLOCK))
	}
	return s
}

pub fn (s TcpSocket) set_option_bool(opt SocketOption, value bool) ? {
	// TODO reenable when this `in` operation works again
	// if opt !in opts_can_set {
	// 	return err_option_not_settable
	// }

	// if opt !in opts_bool {
	// 	return err_option_wrong_type
	// }

	socket_error(C.setsockopt(s.handle, C.SOL_SOCKET, int(opt), &value, sizeof(bool)))?

	return none
}

pub fn (s TcpSocket) set_option_int(opt SocketOption, value int) ? {
	socket_error(C.setsockopt(s.handle, C.SOL_SOCKET, int(opt), &value, sizeof(int)))?

	return none
}

fn (s TcpSocket) close() ? {
	return shutdown(s.handle)
}

fn (s TcpSocket) @select(test Select, timeout time.Duration) ?bool {
	return @select(s.handle, test, timeout)
}

const (
	connect_timeout = 5 * time.second
)

fn (s TcpSocket) connect(a string) ? {
	addr := resolve_addr(a, .inet, .tcp)?
	
	res := C.connect(s.handle, &addr.addr, addr.len)

	if res == 0 {
		return none
	}

	errcode := error_code()

	if errcode == error_ewouldblock {
		write_result := s.@select(.write, connect_timeout)?
		if write_result {
			// succeeded
			return none
		}
		except_result := s.@select(.except, connect_timeout)?
		if except_result {
			return err_connect_failed
		}
		// otherwise we timed out
		return err_connect_timed_out
	}

	wrap_error(errcode)?

	return none
}